
// project.v — TinyTapeout wrapper (top)
`default_nettype none
module tt_um_sfg_cdr (
  input  wire [7:0] ui_in,
  output wire [7:0] uo_out,
  input  wire [7:0] uio_in,
  output wire [7:0] uio_out,
  output wire [7:0] uio_oe,
  input  wire       ena,
  input  wire       clk,      // 50 MHz
  input  wire       rst_n
);
  // ---- your core (unchanged) ----
  wire signed [7:0] y_n = ui_in;
  wire        sample_en;
  wire signed [7:0] x_n;
  wire        d_bb;
  wire [1:0]  d_q2;
  wire signed [15:0] f_n;
  wire signed [31:0] v_ctrl;
  wire signed [31:0] dfcw;

  cdr u_cdr (
    .clk(clk), .rst_n(rst_n), .y_n(y_n),
    .sample_en(sample_en), .x_n(x_n), .d_bb(d_bb), .d_q2(d_q2),
    .f_n(f_n), .v_ctrl(v_ctrl), .dfcw(dfcw)
  );

  // ---- 50% duty recovered clock (toggle on baud strobe) ----
  reg rec_clk;
  always @(posedge clk or negedge rst_n)
    if (!rst_n) rec_clk <= 1'b0;
    else if (sample_en) rec_clk <= ~rec_clk;

  // ---- outputs (quiet when ena=0) ----
  wire [7:0] outs = {
    dfcw[31],     // [7]
    v_ctrl[31],   // [6]
    d_q2[1],      // [5]
    d_q2[0],      // [4]
    d_bb,         // [3]
    x_n[7],       // [2]
    rec_clk,      // [1] REC_CLK 50% duty
    sample_en     // [0] SAMPLE_EN pulse
  };

  assign uo_out  = ena ? outs : 8'h00;
  assign uio_out = 8'h00;
  assign uio_oe  = 8'h00;
endmodule
`default_nettype wire
